`timescale 1ns / 1ps

module Main_Comparator_STRAIT (
    input  wire        clk,
    input  wire        rst,
    input  wire [31:0] accum_out, // RAM �Ǵ� Bus���� ���� ��
    input  wire [31:0] expected,  // ROM���� ���� ����
    output reg         ERROR
);

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            ERROR <= 0;
        end else begin
            // [������ ��] 
            // 1. �����Ͱ� 0�� ���� "���� �����Ͱ� �� �Դ�"�� ���� �����մϴ�.
            // 2. �����Ͱ� 0�� �ƴѵ�(��ȿ�ѵ�) ����(expected)�� �ٸ��� �����Դϴ�.
            // (����: �׽�Ʈ ������ ������ ��� 0�� �ƴ� ������ �����Ǿ� �ֽ��ϴ�)
            if ((accum_out != 32'd0) && (accum_out !== expected)) begin
                ERROR <= 1;
            end
            // �ѹ� ������ ���� 1�� ���� (Sticky)
        end
    end

endmodule