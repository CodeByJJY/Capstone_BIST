`timescale 1ns / 1ps

module tb_System_Top;

    // =========================================================
    // 1. �ùķ��̼� �Ķ���� ����
    // =========================================================
    parameter CLK_PERIOD   = 10; // 100MHz
    parameter ARRAY_SIZE   = 16; 
    parameter NUM_PATTERNS = 16; 
    
    parameter A_WIDTH = 8;
    parameter W_WIDTH = 8;
    parameter P_WIDTH = 32;

    // =========================================================
    // 2. ���� ���� ��ȣ
    // =========================================================
    reg clk;
    reg rst;
    reg start;

    // =========================================================
    // 3. DUT 1: BICS-BIST (����) ��ȣ
    // =========================================================
    wire bics_done;
    wire bics_final_error;
    
    reg  [(ARRAY_SIZE*ARRAY_SIZE)-1:0] bics_pe_disable_bus;
    reg  [(A_WIDTH*ARRAY_SIZE)-1:0]    bics_flat_in_a;
    reg  [(W_WIDTH*ARRAY_SIZE)-1:0]    bics_flat_in_w;
    reg  [(P_WIDTH*ARRAY_SIZE)-1:0]    bics_flat_in_p;
    wire [(A_WIDTH*ARRAY_SIZE)-1:0]    bics_flat_out_a;
    wire [(W_WIDTH*ARRAY_SIZE)-1:0]    bics_flat_out_w;

    // =========================================================
    // 4. DUT 2: STRAIT (����) ��ȣ
    // =========================================================
    wire strait_done;
    // [����] error_count ��Ʈ ���� (���� ��⿡ �����Ƿ�)
    reg  [1:0] strait_bist_mode;

    // =========================================================
    // 5. ���� ���� ����
    // =========================================================
    integer start_time;
    integer bics_end_time;
    integer strait_end_time;
    
    integer bics_cycles;
    integer strait_cycles;

    // =========================================================
    // 6. Ŭ�� ����
    // =========================================================
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end

    // =========================================================
    // 7. DUT �ν��Ͻ�ȭ
    // =========================================================

    // --- [DUT 1] BICS-BIST System ---
    BIST_System_Top_BICS #(
        .ARRAY_SIZE(ARRAY_SIZE),
        .NUM_PATTERNS(NUM_PATTERNS),
        .A_WIDTH(A_WIDTH),
        .W_WIDTH(W_WIDTH),
        .P_WIDTH(P_WIDTH)
    ) dut_bics (
        .clk(clk),
        .rst(rst),
        .start(start),
        .bist_done(bics_done),
        .final_error(bics_final_error),
        .pe_disable_bus(bics_pe_disable_bus),
        .flat_array_in_a(bics_flat_in_a),
        .flat_array_in_w(bics_flat_in_w),
        .flat_array_in_p(bics_flat_in_p),
        .flat_array_out_a(bics_flat_out_a),
        .flat_array_out_w(bics_flat_out_w)
    );

    // --- [DUT 2] STRAIT System ---
    System_Top_STRAIT dut_strait (
        .clk(clk),
        .reset(rst),           
        .bist_en(start),       
        .bist_mode(strait_bist_mode),
        // [����] error_count ���� ���� (�� �κ��� ���� �����̾���)
        .done(strait_done)
    );

    // =========================================================
    // 8. Watchdog (Ÿ�Ӿƿ�)
    // =========================================================
    initial begin
        #(CLK_PERIOD * 5000);
        $display("\n[Time %0t] Simulation Timeout!", $time);
        $finish;
    end

    // =========================================================
    // 9. ���� �׽�Ʈ �ó�����
    // =========================================================
    initial begin
        // --- �ʱ�ȭ ---
        $display("============================================================");
        $display("   BICS vs STRAIT Fairness Benchmark Simulation Start");
        $display("============================================================");

        rst = 1;
        start = 0;
        
        bics_pe_disable_bus = 0;
        bics_flat_in_a = 0;
        bics_flat_in_w = 0;
        bics_flat_in_p = 0;
        strait_bist_mode = 2'b01;

        // --- ���� ���� ---
        #(CLK_PERIOD * 5);
        rst = 0;
        #(CLK_PERIOD * 5);

        // --- �׽�Ʈ ���� ---
        start = 1;
        start_time = $time;
        $display("[Time %0t] Test START!", $time);

        // --- �Ϸ� ��� ---
        fork
            // Thread 1: BICS
            begin
                wait(bics_done);
                bics_end_time = $time;
                bics_cycles = (bics_end_time - start_time) / CLK_PERIOD;
                $display("[Time %0t] BICS-BIST Completed! (Cycles: %0d)", $time, bics_cycles);
            end

            // Thread 2: STRAIT
            begin
                wait(strait_done);
                strait_end_time = $time;
                strait_cycles = (strait_end_time - start_time) / CLK_PERIOD;
                $display("[Time %0t] STRAIT Completed! (Cycles: %0d)", $time, strait_cycles);
            end
        join

        #(CLK_PERIOD * 10);

        // =========================================================
        // 10. ���� ��� ����Ʈ
        // =========================================================
        $display("\n============================================================");
        $display("                  FINAL BENCHMARK REPORT                    ");
        $display("============================================================");
        
        // 1. �ӵ� ��
        $display("1. Test Speed (Latency):");
        $display("   - BICS-BIST : %5d Cycles", bics_cycles);
        $display("   - STRAIT    : %5d Cycles", strait_cycles);
        
        if (bics_cycles < strait_cycles)
            $display("   >> RESULT: BICS is FASTER!");
        else
            $display("   >> RESULT: STRAIT is FASTER (Unexpected?)");

        // 2. ���(����) ��
        $display("\n2. Error Status:");
        
        // BICS ��� Ȯ��
        if (bics_final_error == 0)
            $display("   - BICS Status   : PASS");
        else
            $display("   - BICS Status   : FAIL");

        // STRAIT ��� Ȯ�� (������: ���� ��ȣ ���� ����)
        // dut_strait ������ 'err_flag' ���̾ ���� �о�� (Hierarchical Reference)
        if (dut_strait.err_flag == 0) 
            $display("   - STRAIT Status : PASS (Internal signal checked)");
        else 
            $display("   - STRAIT Status : FAIL (Internal signal checked)");

        $display("============================================================\n");
        $finish;
    end

endmodule